module Task1(a,b,c,d,out);
input wire	a,b,c,d;
output wire	out;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;

assign	SYNTHESIZED_WIRE_1 = ~(c & SYNTHESIZED_WIRE_0);
assign	SYNTHESIZED_WIRE_6 =  ~b;
assign	SYNTHESIZED_WIRE_3 = ~(d | a);
assign	out = ~(SYNTHESIZED_WIRE_1 | SYNTHESIZED_WIRE_2 | SYNTHESIZED_WIRE_3);
assign	SYNTHESIZED_WIRE_4 =  ~a;
assign	SYNTHESIZED_WIRE_5 =  ~c;
assign	SYNTHESIZED_WIRE_2 = ~(b | SYNTHESIZED_WIRE_4 | SYNTHESIZED_WIRE_5);
assign	SYNTHESIZED_WIRE_0 = ~(SYNTHESIZED_WIRE_6 & a);

endmodule
