module Task2(z,y,out);
input wire	z,y;
output wire	out;
assign	out = z & y;
endmodule
