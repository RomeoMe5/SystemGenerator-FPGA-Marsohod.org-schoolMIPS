{% extends "base" %}
{% block body %}
module {{ project_name }}(
);

//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================

endmodule
{% endblock %}
